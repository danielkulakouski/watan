1
5 5 3 5 6 g 1 2 3 4 5 6 7 8 c 4 1
6 5 6 4 5 g 0 10 c 10 1 2 2 6 3
4 11 1 2 2 12
1
